//! Protection Unit package
package pu_pkg;
    typedef struct packed {
        logic read;
        logic write;
    } policy_entry_t;
endpackage
