LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

PACKAGE Common IS
    TYPE READ_WRITE_ENTRY_TYPE IS RECORD
        READ : STD_LOGIC;
        WRITE : STD_LOGIC;
    END RECORD;

    TYPE POLICY_TYPE IS ARRAY (natural range <>, natural range <>) of READ_WRITE_ENTRY_TYPE;
END PACKAGE;

PACKAGE BODY Common IS
END PACKAGE BODY;